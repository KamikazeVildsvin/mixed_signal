// sch_path: /Users/nlv/Documents/DTU/9.Semester/IC-Open-Source/xschem-projects/mixed_signal/mixed_signal
module mixed_signal
(
  output wire Y,
  input wire A1,
  input wire A2,
  input wire B1
);
o21ai_0
x2 ( 
 .A1( A1 ),
 .A2( A2 ),
 .B1( B1 ),
 .Y( Y )
);

endmodule
